`timescale	1ns	/	1ps
module	uart_rx(
	input			clk,														//50MHz主时钟
	input			rst_n,														//低电平复位信号
	input			rs232_rx,													//RS232接收的数据信号
	input			clk_bps,													//此时clk_bps的高电平为接收数据的中间采样点
	output			bps_start,													//接收到信号后，波特率时钟启动信号置位
	output	[7:0]	rx_data,													//接收数据寄存器，保存直到下一个数据来到
	output	reg		rx_int														//接收数据中断信号，接收到数据期间始终为高电平，传送给串口发送模块，
																				//使得串口正在进行数据接收的时候，发送模块不工作，
																				//避免了一个完整数据（1起始位，8数据位，1停止位）还没有完全接收时，
																				//发送模块就已经将不正确的数据传送出去
);

/******************************************************************
*边沿检测程序————检测rs232_rx信号，即串口线上传向FPGA的信号下降沿。
*这个下降沿信号表示一个串口数据帧的开始
*******************************************************************/
	reg				rs232_rx0,rs232_rx1,rs232_rx2,rs232_rx3;					//接收数据寄存器，滤波用
	wire			neg_rs232_rx;												//表示数据线接收到下降沿
	
always	@(posedge	clk	or	negedge	rst_n)
	begin
		if(!rst_n)
			begin
				rs232_rx0	<=	1'b0;
				rs232_rx1	<=	1'b0;
				rs232_rx1	<=	1'b0;
				rs232_rx2	<=	1'b0;
			end
		else
			begin
				rs232_rx0	<=	rs232_rx;
				rs232_rx1	<=	rs232_rx0;
				rs232_rx2	<=	rs232_rx1;
				rs232_rx3	<=	rs232_rx2;
			end
	end
//下面下的降沿检测可以滤掉<20ns~40ns的毛刺（包括高脉冲和低脉冲毛刺），
//在这里就是利用资源来换取稳定（当然我们所需有效低脉冲信号肯定是远远大于40ns的）
assign	neg_rs232_rx	=	rs232_rx3	&	rs232_rx2	&	~rs232_rx1	&	~rs232_rx0	;
//接收到下降沿后neg_rs232_rx置高一个时钟周期

/**************************************************************
*波特率时钟启动信号设置
**************************************************************/
	reg					bps_start_r;
	reg		[3:0]		num;													//移位次数
	// reg					rx_int;													//接收数据中断信号，接收到数据期间始终为高电平

always	@(posedge	clk	or	negedge	rst_n)
	begin
		if(!rst_n)
			begin
				bps_start_r		<=		1'b0;
				rx_int			<=		1'b0;
			end
		else
			if(neg_rs232_rx)													//接收到串口接收线rs232_rx的下降沿标志信号
				begin															
					bps_start_r		<=		1'b1;								//启动串口准备数据接收
					rx_int			<=		1'b1;								//接收数据中断信号使能
				end						
			else						
				if(num	==	4'd12)												//接收完有用数据信息
					begin														
						bps_start_r		<=		1'b0;							//数据接收完毕，释放波特率启动信号
						rx_int			<=		1'b0;							//接收数据终端信号关闭
					end			
	end
assign	bps_start	=	bps_start_r;
/**********************************************************
*数据接模块
***********************************************************/
	reg		[7:0]		rx_data_r;												//串口接收数据寄存器，保存直至下一个数据到来
	reg		[7:0]		rx_temp_data;											//当前接收数据寄存器
	
always	@(posedge	clk	or	negedge	rst_n)
	if(!rst_n)
		begin
			rx_temp_data	<=	8'd0;
			num				<=	4'd0;
			rx_data_r		<=	8'd0;
		end
	else
		begin																	//接收数据处理
			if(clk_bps)
				begin															//读取并保存数据，接收数据为1起始位，8数据位，1或2结束位
					num		<=		num	+	1'b1;
						case(num)
							4'd1:	rx_temp_data[0]		<=		rs232_rx;		//	锁存第0bit
							4'd2:	rx_temp_data[1]		<=		rs232_rx;		//	锁存第1bit
							4'd3:	rx_temp_data[2]		<=		rs232_rx;		//	锁存第2bit
							4'd4:	rx_temp_data[3]		<=		rs232_rx;		//	锁存第3bit
							4'd5:	rx_temp_data[4]		<=		rs232_rx;		//	锁存第4bit
							4'd6:	rx_temp_data[5]		<=		rs232_rx;		//	锁存第5bit
							4'd7:	rx_temp_data[6]		<=		rs232_rx;		//	锁存第6bit
							4'd8:	rx_temp_data[7]		<=		rs232_rx;		//	锁存第7bit
							default: ;
						endcase
				end
			else
				if(num	==	4'd12)
					begin														//我们的标准接收模式下只有1+8+1(2)=11bit的有效数据
						num				<=		4'd0;							//接收到STOP位之后结束，num清零
						rx_data_r		<=		rx_temp_data;					//把锁存的数据送到数据寄存器rx_data中
					end
		end
assign	rx_data		=		rx_data_r;
	
endmodule










