module	speed_select(
	input				clk,
	input				rst_n,
	input				bps_start,			//接收到数据后，波特率时钟启动信号置位，波特率时钟启动信号
	output				clk_bps				//接收或者发送数据位的中间采样点
);

`define		BPS_PARA	5207				//9600波特率时分频计数值
`define		BPS_PARA2	2603				//9600波特率时分频计数值的一半，用于数据采样

	reg		[12:0]		cnt;					//分频计数
	reg					clk_bps_r;				//波特率时钟寄存器

always	@(posedge	clk	or	negedge	rst_n)
	if(!rst_n)
		cnt		<=		13'd0;
	else
		if((cnt	==	`BPS_PARA)	||	!bps_start)
			cnt		<=		13'd0;				
		else
			cnt		<=	cnt		+1'b1;
			
always	@(posedge	clk	or	negedge	rst_n)
	if(!rst_n)
		clk_bps_r	<=	1'b0;
	else
		if(cnt	==	`BPS_PARA2)
			clk_bps_r	<=	1'b1;
		else
			clk_bps_r	<=	1'b0;
			
assign	clk_bps	=	clk_bps_r;

endmodule

/*
parameter         bps9600     = 5207,    //波特率为9600bps
                 bps19200     = 2603,    //波特率为19200bps
                bps38400     = 1301,    //波特率为38400bps
                bps57600     = 867,    //波特率为57600bps
                bps115200    = 433;    //波特率为115200bps 

parameter        bps9600_2     = 2603,
                bps19200_2    = 1301,
                bps38400_2    = 650,
                bps57600_2    = 433,
                bps115200_2 = 216;  
*/